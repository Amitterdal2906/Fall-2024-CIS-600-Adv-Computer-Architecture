library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;  

entity Instruction_Memory is
port (
 pc: in std_logic_vector(31 downto 0);
 im_instruction: out  std_logic_vector(31 downto 0)
);
end Instruction_Memory;

architecture Behavioral of Instruction_Memory is
signal rom_addr: std_logic_vector(31 downto 0);

 type ROM_type is array (0 to 28 ) of std_logic_vector(31 downto 0);
 constant rom_data: ROM_type:=(
--	0 => "10001100001000000000000000000000",  --[lw r0,0(r0)]
--	1 => "10001100001000000000000000000001",  --[lw r0,1(r0)]
--	2 => "10010100000000000000000000000001",  --[lhu r0,1(r0)]
--   3 => "10011100000000000000000000000001",  --[lh  r0,1(r0)]
--	4 => "10010000000000000000000000000000",  --[lbu r0,0(r0)]
--	5 => "10011000000000000000000000000000",  --[lb  r0,0(r0)]
--	6 => "10001100000000000000000000000011",  --[lw r0,3(r0)]
--	7 => "10101100111000000000000000000011",  --[sw r7,3(r0)]
--	8 => "10001100000000000000000000000011",  --[lw r0,3(r0)]
--	9 => "10001100000000000000000000000100",  --[lw r0,4(r0)]
--	10 => "10100100110000000000000000000100", --[sh r6,4(r0)]
--	11 => "10001100000000000000000000000100", --[lw r0,4(r0)]
--	12 => "10001100000000000000000000000101", --[lw r0,5(r0)]
--	13 => "10100000101000000000000000000101", --[sb r5,5(r0)]
--	14 => "10001100000000000000000000000101", --[lw r0,5(r0)]

	
   0 =>  "00000000011000100000000000100000", --[add r3,r2,r0]
   1 =>  "00000000011000100000000000100010", --[sub r3,r2,r0]
   2 =>  "00000000111001100000000000100100", --[and r7,r6,r0]
   3 =>  "00000000101001100000000000100101", --[or r5,r6,r0]
   4 =>  "00000000011000100000000000100110", --[xor r3,r2,r0]
   5 =>  "00000000101000100000000000100111", --[nor r5,r2,r0]
   6 =>  "00000000011000100000000000101010", --[slt r3,r2,r0]
	7 =>  "00000000011011000000000000111011", --[sltu r3,r4,r0]
	8 =>  "00000000011000010000000000000000", --[sll r0,r3,1]
	9 =>  "00000000011000010000000000000010", --[srl r0,r3,1]
	10 => "00000000011000010000000000000011", --[sra r0,r3,1]
	11 => "00000000100000010000000000000111", --[srav r4 1]
	12 => "00000000001000100000000000000100", --[sllv r1 2]
	13 => "00000000100000100000000000000101", --[srlv r4 2]
	14 => "10010100000000000000000000000001", --[lhu r0,1(r0)]
	15 => "10011100000000000000000000000001", --[lh  r0,1(r0)]
	16 => "10010000000000000000000000000000", --[lbu r0,0(r0)]
	17 => "10011000000000000000000000000000", --[lb  r0,0(r0)]	
	18 => "10001100001000000000000000000000", --[lw r0,0(r0)]
	19 => "10101100111000000000000000000011", --[sw r7,3(r0)]
	20 => "10001100000000000000000000000011", --[lw r0,3(r0)]
	21 => "10100100110000000000000000000100", --[sh r6,4(r0)]
	22 => "10001100000000000000000000000100", --[lw r0,4(r0)]
	23 => "10100000101000000000000000000101", --[sb r5,5(r0)]
	24 => "10001100000000000000000000000101", --[lw r0,5(r0)]
	25 =>  "00000000011001000000000000100001", --[addu r3,r4,r0]
   26 =>  "00000000110001000000000000100011", --[subu r6,r4,r0]
   others => x"00000000"

  );
begin


  im_instruction <= rom_data(to_integer(unsigned(pc)));

end Behavioral;